library verilog;
use verilog.vl_types.all;
entity Excesso3TOBCD_vlg_vec_tst is
end Excesso3TOBCD_vlg_vec_tst;
